module SPLITSTREAMER (

);


endmodule
